/*




*/
module win_checker (clk, reset, );
	
endmodule
