///*
//
//
//
//
//*/
//module legality_checker ();
//	input  logic clk, reset;
//	input  logic 
//	
//	output logic enter_output;
//	
//	// Mux... if it's legal, then enter output is whatever enter is
//	// Else, enter output is just 0
//	
//	
//	
//endmodule
