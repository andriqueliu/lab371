///*
//
//
//
//
//*/
//module pctgFSM (clk, reset, address, HEX);
//	input  logic clk, reset;
//	input  integer address;
//	
//	output logic [6:0] HEX;
//	
//	logic  [9:0] pctgReg;
//	
//	percentageDisplay pctgDisplay (.HEX5(HEX), .percent(pctgReg));
//	
//	// 
//	// 
//	always_comb begin
//		case (address)
//			
//		endcase
//	end
//	
//endmodule
