// nios2_tutorial.v

// Generated using ACDS version 14.0 200 at 2017.02.15.15:15:38

`timescale 1 ps / 1 ps
module nios2_tutorial (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule
