/*
EE 371 Lab 2 Project
Andrique Liu, Nikhil Grover, Emraj Sidhu


*/
module inputModule ();

endmodule
