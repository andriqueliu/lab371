// nios2_tutorial.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module nios2_tutorial (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule
